
`ifndef IOB_7KS_V
`define IOB_7KS_V


/**
 * The chip's configurable input/output control blocks
 *
 * MAX7000E and MAX7000S devices
 */
module io_control_block
        (

        ;)

// TODO: see device family datasheet page 15

endmodule

`endif
