
`ifndef EPM7032S_VH
`define EPM7032S_VH

`define LAB_COUNT                       2
`define IO_COUNT                        32

`define BITS_PER_PIA_TO_LAB_ROUTER      4

`endif
