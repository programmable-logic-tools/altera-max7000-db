
`ifndef IOB_7K_V
`define IOB_7K_V


/**
 * The chip's configurable input/output control blocks
 *
 * EPM7032, EPM7064 and EPM7096 devices
 */
module io_control_block
        (

        ;)

// TODO: see device family datasheet page 15

endmodule

`endif
