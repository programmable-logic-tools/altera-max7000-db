
`ifndef MAX7000_FAMILY_VH
`define MAX7000_FAMILY_VH

`endif
