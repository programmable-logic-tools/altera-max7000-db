
`ifndef DEVICE_SPECIFIC_PARAMETERS

`include "epm7032s.vh"

`endif
