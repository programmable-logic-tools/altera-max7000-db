
`ifndef MAX7000_VH
`define MAX7000_VH


`define NUM_GLOBAL_OUTPUT_ENABLE_SIGNALS    6


`endif
