
`ifndef PRIMITIVES_VH
`define PRIMITIVES_VH

`include "iob.v"
`include "lab.v"
`include "macrocell.v"
`include "pia_router.v"
`include "pia.v"
`include "product_term.v"

`endif
